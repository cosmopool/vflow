module commands
