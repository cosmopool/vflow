module commands

pub struct ModuleProperties {
	command string
	options []string
	flags   []string
	usage   string
}
