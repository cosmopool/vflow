module vflow


fn test_check_requirements(){
  /* assert vflow.check_requirements() == true */
  assert true == true
}
